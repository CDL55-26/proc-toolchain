module Bit_OR(
    output [31:0] Or_out,
    input [31:0] A,
    input [31:0] B
);

or or_0(Or_out[0],A[0],B[0]);
or or_1(Or_out[1],A[1],B[1]);
or or_2(Or_out[2],A[2],B[2]);
or or_3(Or_out[3],A[3],B[3]);
or or_4(Or_out[4],A[4],B[4]);
or or_5(Or_out[5],A[5],B[5]);
or or_6(Or_out[6],A[6],B[6]);
or or_7(Or_out[7],A[7],B[7]);
or or_8(Or_out[8],A[8],B[8]);
or or_9(Or_out[9],A[9],B[9]);
or or_10(Or_out[10],A[10],B[10]);
or or_11(Or_out[11],A[11],B[11]);
or or_12(Or_out[12],A[12],B[12]);
or or_13(Or_out[13],A[13],B[13]);
or or_14(Or_out[14],A[14],B[14]);
or or_15(Or_out[15],A[15],B[15]);
or or_16(Or_out[16],A[16],B[16]);
or or_17(Or_out[17],A[17],B[17]);
or or_18(Or_out[18],A[18],B[18]);
or or_19(Or_out[19],A[19],B[19]);
or or_20(Or_out[20],A[20],B[20]);
or or_21(Or_out[21],A[21],B[21]);
or or_22(Or_out[22],A[22],B[22]);
or or_23(Or_out[23],A[23],B[23]);
or or_24(Or_out[24],A[24],B[24]);
or or_25(Or_out[25],A[25],B[25]);
or or_26(Or_out[26],A[26],B[26]);
or or_27(Or_out[27],A[27],B[27]);
or or_28(Or_out[28],A[28],B[28]);
or or_29(Or_out[29],A[29],B[29]);
or or_30(Or_out[30],A[30],B[30]);
or or_31(Or_out[31],A[31],B[31]);

endmodule